//=====================================================================
// Project: 4 core MESI cache design
// File Name: test_lib.svh
// Description: Base test class and list of tests
// Designers: Venky & Suru
//=====================================================================
//TODO: add your testcase files in here
`include "base_test.sv"
`include "read_miss_icache.sv"
`include "read_hit_icache.sv"
`include "read_miss_dcache.sv"
`include "read_hit_dcache.sv"
`include "write_miss_dcache.sv"
`include "write_hit_dcache.sv"
